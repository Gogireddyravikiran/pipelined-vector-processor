`timescale 1 ns / 1 ps

module testbench;
	reg clk =1 ;
	reg reset ;
    always #5 clk = ~clk;
    reg [7:0] instruction;
    reg alu_enb;
    wire alu_done;

    reg [511:0] opA;
    reg [511:0] opB;
    reg [511:0] opC;
    wire [511:0] alu_out;

    reg [31:0] SEW;
    reg [3:0] vap;
    reg [31:0] vlmax;
    
   vector_alu dut(clk, reset, instruction,alu_enb,alu_done,opA,opB,opC,alu_out,SEW,vap,vlmax);


    localparam instr_vadd__vv = 8'h00 ;
    localparam instr_vsub__vv = 8'h01 ;
    localparam instr_vmul__vv = 8'h02 ;
    localparam instr_vmacc_vv = 8'h03 ;
    localparam instr_vmulvarp = 8'h04 ;
    localparam instr_vaddvarp = 8'h05 ;
    localparam instr_vsubvarp = 8'h06 ;
    localparam instr_vmaccvarp = 8'h07 ; 



    initial begin
        
        reset = 1;
        #(10);
        reset = 0;
       // opA         = 512'b00001000110010100111010000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        //opB         = 512'b00001000110010100111010000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        //opC         = 512'b00001000110010100111010000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

        //opB         = 512'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010100000101010001;
        //opC         = 512'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010001010100000100;
//       opA={{480{1'b0}},32'h87654321} ;
//       opB={{480{1'b0}},32'h11111111} ;
//       opC={{480{1'b0}},32'h00000000} ;

         opB = {32'h87654321,480'd0};
         opA = {128'h11111111111111111111111111111111,384'd0};
         opC = 512'd0;
       
        instruction = instr_vmacc_vv;
 
        alu_enb = 1;
        SEW         = 16;
        vap         = 3;
     
       
        #(350);

        $finish;
    end


endmodule